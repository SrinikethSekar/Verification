interface flipflop;
  
  logic clk;
  logic rst;
  logic data;
  logic q_b;
  logic q;
  
endinterface

  
